lpm_dff1_inst : lpm_dff1 PORT MAP (
		aclr	 => aclr_sig,
		aload	 => aload_sig,
		aset	 => aset_sig,
		clock	 => clock_sig,
		data	 => data_sig,
		enable	 => enable_sig,
		q	 => q_sig
	);
