lpm_dff0_inst : lpm_dff0 PORT MAP (
		aclr	 => aclr_sig,
		clock	 => clock_sig,
		data	 => data_sig,
		enable	 => enable_sig,
		sclr	 => sclr_sig,
		q	 => q_sig
	);
